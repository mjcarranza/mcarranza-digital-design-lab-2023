
module CompuertaAND #(parameter N=2) (
  input wire [N-1:0] a, // Entradas de la compuerta AND
  output wire out       // Salida de la compuerta AND
);

  assign out = &a; // La salida es la operación AND de todas las entradas a través de la función "&".

endmodule