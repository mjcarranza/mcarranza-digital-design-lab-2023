module BuscaMinas();
	
	



endmodule
